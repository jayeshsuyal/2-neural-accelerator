`ifndef NEURAL_BASE_SEQ_SV
`define NEURAL_BASE_SEQ_SV

class neural_base_seq extends uvm_sequence #(neural_tx);
    `uvm_object_utils(neural_base_seq)



endclass
`endif